`include "addr_intf.sv"
`include "addr_dut.sv"
`include "addr_trans.sv"
`include "addr_sequence1.sv"
`include "addr_driver.sv"
`include "addr_monitor1.sv"
`include "addr_agent1.sv"
`include "addr_env.sv"
`include "addr_test.sv"
